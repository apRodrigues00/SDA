library IEEE;
use IEEE.std_logic_1164.all;

entity decoder is
port(
	enable		:  in std_logic;
	sel			:	in std_logic_vector(4 downto 0);
	write_reg	:	out std_logic_vector(31 downto 0)
	);
end entity;

architecture arc_decoder of decoder is

begin
	process(enable, sel)
	begin

	 if enable='1' then 
		case sel is  
			when "00000" => write_reg <= "00000000000000000000000000000001" ;
			when "00001" => write_reg <= "00000000000000000000000000000010" ;
			when "00010" => write_reg <= "00000000000000000000000000000100" ;
			when "00011" => write_reg <= "00000000000000000000000000001000" ;
			when "00100" => write_reg <= "00000000000000000000000000010000" ;
			when "00101" => write_reg <= "00000000000000000000000000100000" ;
			when "00110" => write_reg <= "00000000000000000000000001000000" ;
			when "00111" => write_reg <= "00000000000000000000000010000000" ;
			when "01000" => write_reg <= "00000000000000000000000100000000" ;
			when "01001" => write_reg <= "00000000000000000000001000000000" ;
			when "01010" => write_reg <= "00000000000000000000010000000000" ;
			when "01011" => write_reg <= "00000000000000000000100000000000" ;
			when "01100" => write_reg <= "00000000000000000001000000000000" ;
			when "01101" => write_reg <= "00000000000000000010000000000000" ;
			when "01110" => write_reg <= "00000000000000000100000000000000" ;
			when "01111" => write_reg <= "00000000000000001000000000000000" ;
			when "10000" => write_reg <= "00000000000000010000000000000000" ;
			when "10001" => write_reg <= "00000000000000100000000000000000" ;
			when "10010" => write_reg <= "00000000000001000000000000000000" ;
			when "10011" => write_reg <= "00000000000010000000000000000000" ;
			when "10100" => write_reg <= "00000000000100000000000000000000" ;
			when "10101" => write_reg <= "00000000001000000000000000000000" ;
			when "10110" => write_reg <= "00000000010000000000000000000000" ;
			when "10111" => write_reg <= "00000000100000000000000000000000" ;
			when "11000" => write_reg <= "00000001000000000000000000000000" ;
			when "11001" => write_reg <= "00000010000000000000000000000000" ;
			when "11010" => write_reg <= "00000100000000000000000000000000" ;
			when "11011" => write_reg <= "00001000000000000000000000000000" ;
			when "11100" => write_reg <= "00010000000000000000000000000000" ;
			when "11101" => write_reg <= "00100000000000000000000000000000" ;
			when "11110" => write_reg <= "01000000000000000000000000000000" ;
			when "11111" => write_reg <= "10000000000000000000000000000000" ;
		end case;
		else 
			write_reg <= "00000000000000000000000000000000";
		end if;
	end process;
end architecture;