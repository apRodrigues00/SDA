library verilog;
use verilog.vl_types.all;
entity somador_nbits_vlg_vec_tst is
end somador_nbits_vlg_vec_tst;
